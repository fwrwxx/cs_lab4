module Ex2_OR(x1,x2,f);
input x1,x2;
output f;
assign f = ( x1 & ~x2 )|( ~x1 & x2 );
endmodule

module Ex2_OR(x1,x2,x3,f);
  input x1,x2,x3;
  output f;
  wire f;
  assign f = ( ~x3 & ~x2 )|( x1 & ( x3 ^ x2) );
endmodule

module Ex2_OR(x1,x2,x3,f);
  input x1,x2,x3;
  output f;
  wire f;
  assign f = ( ~x1 )&( x2 | x3);
endmodule
